* Extracted by KLayout with SG13G2 LVS runset on : 08/05/2024 12:11

* cell IDSM2_t1_inner
* pin sub!
.SUBCKT IDSM2_t1_inner sub!
* device instance $1 r0 *1 85.1,-27.161 sg13_lv_nmos
M$1 sub! \$6 \$3 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $2 r0 *1 80.056,-23.537 sg13_lv_nmos
M$2 \$5 \$6 \$201 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $3 r0 *1 80.057,-18.777 sg13_lv_nmos
M$3 sub! \$198 \$16 sub! sg13_lv_nmos W=1.9999999999999996 L=0.9999999999999998
* device instance $4 r0 *1 82.656,-18.777 sg13_lv_nmos
M$4 sub! \$5 \$17 sub! sg13_lv_nmos W=1.9999999999999996 L=0.9999999999999998
* device instance $5 r0 *1 106.28,-17.578 sg13_lv_nmos
M$5 \$31 \$88 \$68 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $6 r0 *1 106.59,-17.578 sg13_lv_nmos
M$6 \$68 \$18 sub! sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $7 r0 *1 107.17,-17.193 sg13_lv_nmos
M$7 sub! \$81 \$32 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $8 r0 *1 115.01,-17.578 sg13_lv_nmos
M$8 \$34 \$35 sub! sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $9 r0 *1 115.52,-17.578 sg13_lv_nmos
M$9 sub! \$18 \$58 sub! sg13_lv_nmos W=0.41999999999999993 L=0.12999999999999995
* device instance $10 r0 *1 115.83,-17.578 sg13_lv_nmos
M$10 \$58 \$49 \$35 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $11 r0 *1 117.87,-17.468 sg13_lv_nmos
M$11 sub! \$49 \$37 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $12 r0 *1 116.85,-17.418 sg13_lv_nmos
M$12 sub! \$49 \$36 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $14 r0 *1 118.89,-17.418 sg13_lv_nmos
M$14 sub! \$37 \$38 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $16 r0 *1 80.056,-17.244 sg13_lv_nmos
M$16 \$16 \$30 \$43 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $17 r0 *1 82.656,-17.248 sg13_lv_nmos
M$17 \$17 \$30 \$44 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $18 r0 *1 89.915,-17.364 sg13_lv_nmos
M$18 sub! \$86 \$45 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $19 r0 *1 92.727,-17.39 sg13_lv_nmos
M$19 sub! \$92 \$46 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $20 r0 *1 105.025,-17.398 sg13_lv_nmos
M$20 sub! \$14 \$18 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $21 r0 *1 108.26,-17.513 sg13_lv_nmos
M$21 sub! \$18 \$64 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $22 r0 *1 108.57,-17.513 sg13_lv_nmos
M$22 \$64 \$32 \$47 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $23 r0 *1 111.115,-17.313 sg13_lv_nmos
M$23 sub! \$33 \$48 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $24 r0 *1 112.215,-17.313 sg13_lv_nmos
M$24 sub! \$6 \$33 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $25 r0 *1 113.425,-17.193 sg13_lv_nmos
M$25 \$49 \$33 \$34 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $26 r0 *1 113.96,-17.353 sg13_lv_nmos
M$26 \$32 \$48 \$49 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $27 r0 *1 43.29,-15.84 sg13_lv_nmos
M$27 sub! \$21 \$22 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $31 r0 *1 46.17,-15.84 sg13_lv_nmos
M$31 sub! \$22 \$23 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $35 r0 *1 49.05,-15.84 sg13_lv_nmos
M$35 sub! \$23 \$24 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $39 r0 *1 51.93,-15.84 sg13_lv_nmos
M$39 sub! \$24 \$25 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $43 r0 *1 54.81,-15.84 sg13_lv_nmos
M$43 sub! \$25 \$26 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $47 r0 *1 57.69,-15.84 sg13_lv_nmos
M$47 sub! \$26 \$27 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $51 r0 *1 63.45,-15.84 sg13_lv_nmos
M$51 sub! \$28 \$29 sub! sg13_lv_nmos W=2.9599999999999995 L=0.12999999999999995
* device instance $55 r0 *1 66.27,-15.84 sg13_lv_nmos
M$55 sub! \$29 \$30 sub! sg13_lv_nmos W=5.92 L=0.12999999999999995
* device instance $63 r0 *1 79.854,-16.171 sg13_lv_nmos
M$63 \$43 \$86 \$92 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $64 r0 *1 82.66,-16.155 sg13_lv_nmos
M$64 \$44 \$92 \$86 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $65 r0 *1 89.899,-16.321 sg13_lv_nmos
M$65 \$45 \$88 \$87 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $66 r0 *1 92.728,-16.32 sg13_lv_nmos
M$66 \$46 \$87 \$88 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $67 r0 *1 99.177,-16.341 sg13_lv_nmos
M$67 sub! \$88 \$79 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $68 r0 *1 99.687,-16.391 sg13_lv_nmos
M$68 sub! \$79 \$80 sub! sg13_lv_nmos W=1.4799999999999998 L=0.12999999999999995
* device instance $70 r0 *1 109.345,-16.788 sg13_lv_nmos
M$70 \$31 \$33 \$81 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $71 r0 *1 109.855,-16.788 sg13_lv_nmos
M$71 \$81 \$48 \$47 sub! sg13_lv_nmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $72 r0 *1 36.59,-13.5 sg13_lv_nmos
M$72 sub! \$138 \$78 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $74 r0 *1 38.51,-13.5 sg13_lv_nmos
M$74 sub! \$78 \$127 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $76 r0 *1 40.375,-13.525 sg13_lv_nmos
M$76 \$128 \$127 \$129 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $78 r0 *1 41.405,-13.525 sg13_lv_nmos
M$78 \$128 \$27 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $80 r0 *1 40.375,-15.815 sg13_lv_nmos
M$80 \$84 \$42 \$21 sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $82 r0 *1 41.405,-15.815 sg13_lv_nmos
M$82 \$84 \$78 sub! sub! sg13_lv_nmos W=1.4399999999999997 L=0.12999999999999998
* device instance $84 r0 *1 43.29,-13.5 sg13_lv_nmos
M$84 sub! \$129 \$130 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $88 r0 *1 46.17,-13.5 sg13_lv_nmos
M$88 sub! \$130 \$131 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $92 r0 *1 49.05,-13.5 sg13_lv_nmos
M$92 sub! \$131 \$132 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $96 r0 *1 51.93,-13.5 sg13_lv_nmos
M$96 sub! \$132 \$133 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $100 r0 *1 54.81,-13.5 sg13_lv_nmos
M$100 sub! \$133 \$134 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $104 r0 *1 57.69,-13.5 sg13_lv_nmos
M$104 sub! \$134 \$42 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $108 r0 *1 60.645,-13.525 sg13_lv_nmos
M$108 \$135 \$42 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $110 r0 *1 61.675,-13.525 sg13_lv_nmos
M$110 \$135 \$133 \$139 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $112 r0 *1 60.645,-15.815 sg13_lv_nmos
M$112 \$85 \$27 sub! sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $114 r0 *1 61.675,-15.815 sg13_lv_nmos
M$114 \$85 \$25 \$28 sub! sg13_lv_nmos W=1.4399999999999997
+ L=0.12999999999999998
* device instance $116 r0 *1 63.45,-13.5 sg13_lv_nmos
M$116 sub! \$139 \$136 sub! sg13_lv_nmos W=2.9599999999999995
+ L=0.12999999999999995
* device instance $120 r0 *1 66.27,-13.5 sg13_lv_nmos
M$120 sub! \$136 \$6 sub! sg13_lv_nmos W=5.92 L=0.12999999999999995
* device instance $128 r0 *1 38.045,2.297 sg13_lv_nmos
M$128 sub! \$6 \$188 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $129 r0 *1 39.13,2.397 sg13_lv_nmos
M$129 sub! \$38 \$202 sub! sg13_lv_nmos W=0.5499999999999999
+ L=0.12999999999999995
* device instance $130 r0 *1 39.98,2.302 sg13_lv_nmos
M$130 sub! \$30 \$210 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $131 r0 *1 40.29,2.302 sg13_lv_nmos
M$131 \$210 \$202 \$189 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $132 r0 *1 41.605,2.467 sg13_lv_nmos
M$132 \$203 \$30 \$212 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $133 r0 *1 42.115,2.467 sg13_lv_nmos
M$133 sub! \$38 \$212 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $134 r0 *1 42.625,2.417 sg13_lv_nmos
M$134 sub! \$203 \$190 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $135 r0 *1 47.434,6.03 sg13_lv_nmos
M$135 \$230 \$190 \$236 sub! sg13_lv_nmos W=0.4999999999999999
+ L=0.12999999999999998
* device instance $136 r0 *1 49.852,6.092 sg13_lv_nmos
M$136 \$236 \$6 \$237 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $137 r0 *1 55.875,5.647 sg13_lv_nmos
M$137 sub! \$191 \$191 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $138 r0 *1 55.531,2.757 sg13_lv_nmos
M$138 \$191 \$134 \$204 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $139 r0 *1 56.04,2.757 sg13_lv_nmos
M$139 \$204 \$30 \$192 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $140 r0 *1 60.25,5.632 sg13_lv_nmos
M$140 sub! \$193 \$194 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $141 r0 *1 59.931,2.737 sg13_lv_nmos
M$141 \$193 \$6 \$192 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $142 r0 *1 60.44,2.737 sg13_lv_nmos
M$142 \$192 \$14 \$194 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $143 r0 *1 67.127,2.297 sg13_lv_nmos
M$143 sub! \$30 \$195 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $144 r0 *1 68.212,2.397 sg13_lv_nmos
M$144 sub! \$80 \$205 sub! sg13_lv_nmos W=0.5499999999999999
+ L=0.12999999999999995
* device instance $145 r0 *1 69.062,2.302 sg13_lv_nmos
M$145 sub! \$6 \$215 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $146 r0 *1 69.372,2.302 sg13_lv_nmos
M$146 \$215 \$205 \$196 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $147 r0 *1 70.687,2.467 sg13_lv_nmos
M$147 \$206 \$6 \$214 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $148 r0 *1 71.197,2.467 sg13_lv_nmos
M$148 sub! \$80 \$214 sub! sg13_lv_nmos W=0.6399999999999999
+ L=0.12999999999999995
* device instance $149 r0 *1 71.707,2.417 sg13_lv_nmos
M$149 sub! \$206 \$197 sub! sg13_lv_nmos W=0.7399999999999999
+ L=0.12999999999999995
* device instance $150 r0 *1 76.516,6.03 sg13_lv_nmos
M$150 \$230 \$197 \$231 sub! sg13_lv_nmos W=0.4999999999999999
+ L=0.12999999999999998
* device instance $151 r0 *1 78.934,6.092 sg13_lv_nmos
M$151 \$231 \$30 \$194 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $152 r0 *1 84.957,5.647 sg13_lv_nmos
M$152 sub! \$198 \$198 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $153 r0 *1 84.613,2.757 sg13_lv_nmos
M$153 \$198 \$26 \$207 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $154 r0 *1 85.122,2.757 sg13_lv_nmos
M$154 \$207 \$6 \$199 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $155 r0 *1 89.332,5.632 sg13_lv_nmos
M$155 sub! \$200 \$201 sub! sg13_lv_nmos W=2.4999999999999996
+ L=1.4999999999999996
* device instance $156 r0 *1 89.013,2.737 sg13_lv_nmos
M$156 \$200 \$30 \$199 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $157 r0 *1 89.522,2.737 sg13_lv_nmos
M$157 \$199 \$14 \$201 sub! sg13_lv_nmos W=1.9999999999999996
+ L=0.12999999999999998
* device instance $158 r0 *1 117.585,-12.41 sg13_lv_nmos
M$158 sub! \$38 \$165 sub! sg13_lv_nmos W=1.4799999999999998
+ L=0.12999999999999995
* device instance $160 r0 *1 80.045,-26.542 sg13_lv_pmos
M$160 \$5 \$3 \$201 \$11 sg13_lv_pmos W=5.999999999999998 L=0.12999999999999998
* device instance $163 r0 *1 85.11,-25.486 sg13_lv_pmos
M$163 \$164 \$6 \$3 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $164 r0 *1 40.375,-17.5 sg13_lv_pmos
M$164 \$164 \$42 \$21 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $166 r0 *1 41.405,-17.5 sg13_lv_pmos
M$166 \$164 \$78 \$21 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $168 r0 *1 43.29,-17.5 sg13_lv_pmos
M$168 \$164 \$21 \$22 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $172 r0 *1 46.17,-17.5 sg13_lv_pmos
M$172 \$164 \$22 \$23 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $176 r0 *1 49.05,-17.5 sg13_lv_pmos
M$176 \$164 \$23 \$24 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $180 r0 *1 51.93,-17.5 sg13_lv_pmos
M$180 \$164 \$24 \$25 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $184 r0 *1 54.81,-17.5 sg13_lv_pmos
M$184 \$164 \$25 \$26 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $188 r0 *1 57.69,-17.5 sg13_lv_pmos
M$188 \$164 \$26 \$27 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $192 r0 *1 60.645,-17.5 sg13_lv_pmos
M$192 \$164 \$27 \$28 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $194 r0 *1 61.675,-17.5 sg13_lv_pmos
M$194 \$164 \$25 \$28 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $196 r0 *1 63.45,-17.5 sg13_lv_pmos
M$196 \$164 \$28 \$29 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $200 r0 *1 66.27,-17.5 sg13_lv_pmos
M$200 \$164 \$29 \$30 \$164 sg13_lv_pmos W=8.959999999999999
+ L=0.12999999999999995
* device instance $208 r0 *1 36.58,-11.84 sg13_lv_pmos
M$208 \$164 \$138 \$78 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $210 r0 *1 38.5,-11.84 sg13_lv_pmos
M$210 \$164 \$78 \$127 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $212 r0 *1 40.375,-11.84 sg13_lv_pmos
M$212 \$164 \$127 \$129 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $214 r0 *1 41.405,-11.84 sg13_lv_pmos
M$214 \$164 \$27 \$129 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $216 r0 *1 43.29,-11.84 sg13_lv_pmos
M$216 \$164 \$129 \$130 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $220 r0 *1 46.17,-11.84 sg13_lv_pmos
M$220 \$164 \$130 \$131 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $224 r0 *1 49.05,-11.84 sg13_lv_pmos
M$224 \$164 \$131 \$132 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $228 r0 *1 51.93,-11.84 sg13_lv_pmos
M$228 \$164 \$132 \$133 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $232 r0 *1 54.81,-11.84 sg13_lv_pmos
M$232 \$164 \$133 \$134 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $236 r0 *1 57.69,-11.84 sg13_lv_pmos
M$236 \$164 \$134 \$42 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $240 r0 *1 60.645,-11.84 sg13_lv_pmos
M$240 \$164 \$42 \$139 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $242 r0 *1 61.675,-11.84 sg13_lv_pmos
M$242 \$164 \$133 \$139 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $244 r0 *1 63.45,-11.84 sg13_lv_pmos
M$244 \$164 \$139 \$136 \$164 sg13_lv_pmos W=4.4799999999999995
+ L=0.12999999999999995
* device instance $248 r0 *1 66.27,-11.84 sg13_lv_pmos
M$248 \$164 \$136 \$6 \$164 sg13_lv_pmos W=8.959999999999999
+ L=0.12999999999999995
* device instance $256 r0 *1 78.866,-13.253 sg13_lv_pmos
M$256 \$92 \$30 \$247 \$157 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $257 r0 *1 78.866,-14.683 sg13_lv_pmos
M$257 \$92 \$86 \$247 \$157 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $258 r0 *1 83.665,-13.253 sg13_lv_pmos
M$258 \$86 \$92 \$247 \$183 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $259 r0 *1 83.665,-14.683 sg13_lv_pmos
M$259 \$86 \$30 \$247 \$183 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $260 r0 *1 88.763,-13.253 sg13_lv_pmos
M$260 \$87 \$86 \$164 \$183 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $261 r0 *1 88.763,-14.683 sg13_lv_pmos
M$261 \$87 \$88 \$164 \$183 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $262 r0 *1 93.787,-13.265 sg13_lv_pmos
M$262 \$88 \$87 \$164 \$145 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $263 r0 *1 93.787,-14.695 sg13_lv_pmos
M$263 \$88 \$92 \$164 \$145 sg13_lv_pmos W=3.999999999999999
+ L=0.12999999999999998
* device instance $264 r0 *1 99.177,-14.716 sg13_lv_pmos
M$264 \$164 \$88 \$79 \$164 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $265 r0 *1 99.687,-14.731 sg13_lv_pmos
M$265 \$164 \$79 \$80 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $267 r0 *1 105.035,-15.723 sg13_lv_pmos
M$267 \$164 \$14 \$18 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $268 r0 *1 106.17,-15.988 sg13_lv_pmos
M$268 \$164 \$88 \$31 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $269 r0 *1 106.68,-15.988 sg13_lv_pmos
M$269 \$164 \$18 \$31 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $270 r0 *1 107.13,-15.698 sg13_lv_pmos
M$270 \$164 \$81 \$32 \$164 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $271 r0 *1 108.18,-15.623 sg13_lv_pmos
M$271 \$81 \$18 \$164 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $272 r0 *1 108.915,-15.623 sg13_lv_pmos
M$272 \$164 \$32 \$106 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $273 r0 *1 109.305,-15.623 sg13_lv_pmos
M$273 \$106 \$33 \$81 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $274 r0 *1 109.815,-15.623 sg13_lv_pmos
M$274 \$81 \$48 \$31 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $275 r0 *1 111.515,-15.748 sg13_lv_pmos
M$275 \$48 \$33 \$164 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $276 r0 *1 112.24,-15.748 sg13_lv_pmos
M$276 \$164 \$6 \$33 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $277 r0 *1 114.37,-16.003 sg13_lv_pmos
M$277 \$49 \$48 \$100 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $278 r0 *1 114.75,-16.003 sg13_lv_pmos
M$278 \$100 \$35 \$164 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $279 r0 *1 115.36,-16.003 sg13_lv_pmos
M$279 \$164 \$18 \$35 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $280 r0 *1 115.87,-16.003 sg13_lv_pmos
M$280 \$164 \$49 \$35 \$164 sg13_lv_pmos W=0.41999999999999993
+ L=0.12999999999999995
* device instance $281 r0 *1 117.43,-15.898 sg13_lv_pmos
M$281 \$164 \$49 \$37 \$164 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $282 r0 *1 116.41,-15.838 sg13_lv_pmos
M$282 \$164 \$49 \$36 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $284 r0 *1 113.675,-15.713 sg13_lv_pmos
M$284 \$32 \$33 \$49 \$164 sg13_lv_pmos W=0.9999999999999998
+ L=0.12999999999999998
* device instance $285 r0 *1 118.515,-15.738 sg13_lv_pmos
M$285 \$164 \$37 \$38 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $287 r0 *1 38.055,3.972 sg13_lv_pmos
M$287 \$164 \$6 \$188 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $288 r0 *1 39.13,3.822 sg13_lv_pmos
M$288 \$202 \$38 \$164 \$164 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $289 r0 *1 39.67,3.962 sg13_lv_pmos
M$289 \$164 \$30 \$189 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $290 r0 *1 40.18,3.962 sg13_lv_pmos
M$290 \$189 \$202 \$164 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $291 r0 *1 41.605,4.107 sg13_lv_pmos
M$291 \$164 \$30 \$203 \$164 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $292 r0 *1 42.115,4.107 sg13_lv_pmos
M$292 \$164 \$38 \$203 \$164 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $293 r0 *1 42.625,3.967 sg13_lv_pmos
M$293 \$164 \$203 \$190 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $294 r0 *1 47.838,8.924 sg13_lv_pmos
M$294 \$236 \$188 \$237 \$247 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $297 r0 *1 50.505,9.567 sg13_lv_pmos
M$297 \$236 \$189 \$246 \$247 sg13_lv_pmos W=1.4999999999999998
+ L=0.12999999999999995
* device instance $298 r0 *1 55.886,8.657 sg13_lv_pmos
M$298 \$191 \$191 \$247 \$247 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $302 r0 *1 60.256,8.642 sg13_lv_pmos
M$302 \$194 \$193 \$247 \$247 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $306 r0 *1 67.137,3.972 sg13_lv_pmos
M$306 \$164 \$30 \$195 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $307 r0 *1 68.212,3.822 sg13_lv_pmos
M$307 \$205 \$80 \$164 \$164 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $308 r0 *1 68.752,3.962 sg13_lv_pmos
M$308 \$164 \$6 \$196 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $309 r0 *1 69.262,3.962 sg13_lv_pmos
M$309 \$196 \$205 \$164 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $310 r0 *1 70.687,4.107 sg13_lv_pmos
M$310 \$164 \$6 \$206 \$164 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $311 r0 *1 71.197,4.107 sg13_lv_pmos
M$311 \$164 \$80 \$206 \$164 sg13_lv_pmos W=0.8399999999999999
+ L=0.12999999999999995
* device instance $312 r0 *1 71.707,3.967 sg13_lv_pmos
M$312 \$164 \$206 \$197 \$164 sg13_lv_pmos W=1.1199999999999999
+ L=0.12999999999999995
* device instance $313 r0 *1 76.92,8.924 sg13_lv_pmos
M$313 \$231 \$195 \$194 \$247 sg13_lv_pmos W=5.999999999999998
+ L=0.12999999999999998
* device instance $316 r0 *1 79.587,9.567 sg13_lv_pmos
M$316 \$231 \$196 \$246 \$247 sg13_lv_pmos W=1.4999999999999998
+ L=0.12999999999999995
* device instance $317 r0 *1 84.968,8.657 sg13_lv_pmos
M$317 \$198 \$198 \$247 \$247 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $321 r0 *1 89.338,8.642 sg13_lv_pmos
M$321 \$201 \$200 \$247 \$247 sg13_lv_pmos W=9.999999999999998
+ L=1.4999999999999996
* device instance $325 r0 *1 117.575,-10.75 sg13_lv_pmos
M$325 \$164 \$38 \$165 \$164 sg13_lv_pmos W=2.2399999999999998
+ L=0.12999999999999995
* device instance $327 r0 *1 86.178,-29.692 cap_cmim
C$327 \$5 sub! cap_cmim w=5.77 l=5.77 m=1
* device instance $328 r0 *1 37.283,6.963 cap_cmim
C$328 \$204 \$236 cap_cmim w=5.77 l=5.77 m=1
* device instance $329 r0 *1 66.365,6.963 cap_cmim
C$329 \$207 \$231 cap_cmim w=5.77 l=5.77 m=1
* device instance $330 r0 *1 36.035,14.656 cap_cmim
C$330 \$193 \$204 cap_cmim w=8.16 l=8.16 m=1
* device instance $331 r0 *1 65.117,14.656 cap_cmim
C$331 \$200 \$207 cap_cmim w=8.16 l=8.16 m=1
* device instance $332 r0 *1 52.385,15.898 cap_cmim
C$332 \$192 \$194 cap_cmim w=8.16 l=8.16 m=1
* device instance $333 r0 *1 81.467,15.898 cap_cmim
C$333 \$199 \$201 cap_cmim w=8.16 l=8.16 m=1
.ENDS IDSM2_t1_inner
