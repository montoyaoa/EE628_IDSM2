* Extracted by KLayout with SG13G2 LVS runset on : 30/04/2024 22:43

* cell clock_gen
.SUBCKT clock_gen
.ENDS clock_gen
