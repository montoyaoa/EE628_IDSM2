* Extracted by KLayout with SG13G2 LVS runset on : 05/05/2024 22:53

* cell stage_t1
* pin sub!
.SUBCKT stage_t1 sub!
* device instance $1 r0 *1 12.911,0.09 sg13_lv_nmos
M$1 \$10 \$27 \$18 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $2 r0 *1 13.42,0.09 sg13_lv_nmos
M$2 \$18 \$28 \$11 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $3 r0 *1 8.511,0.11 sg13_lv_nmos
M$3 \$9 \$24 \$17 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $4 r0 *1 9.02,0.11 sg13_lv_nmos
M$4 \$17 \$25 \$18 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $5 r0 *1 13.23,2.985 sg13_lv_nmos
M$5 sub! \$10 \$11 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $6 r0 *1 8.855,3 sg13_lv_nmos
M$6 sub! \$9 \$42 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $7 r0 *1 0.414,3.383 sg13_lv_nmos
M$7 \$35 \$16 \$38 sub! sg13_lv_nmos W=0.4999999999999999 L=0.12999999999999998
* device instance $8 r0 *1 2.832,3.445 sg13_lv_nmos
M$8 \$41 \$5 \$39 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $9 r0 *1 13.236,5.995 sg13_lv_pmos
M$9 \$46 \$10 \$48 \$48 sg13_lv_pmos W=2.4999999999999996 L=1.4999999999999996
* device instance $10 r0 *1 13.236,7.875 sg13_lv_pmos
M$10 \$48 \$10 \$11 \$48 sg13_lv_pmos W=7.499999999999998 L=1.4999999999999996
* device instance $13 r0 *1 8.866,6.01 sg13_lv_pmos
M$13 \$42 \$9 \$48 \$48 sg13_lv_pmos W=9.999999999999998 L=1.4999999999999996
* device instance $17 r0 *1 0.818,6.277 sg13_lv_pmos
M$17 \$41 \$12 \$39 \$48 sg13_lv_pmos W=5.999999999999998 L=0.12999999999999998
* device instance $20 r0 *1 3.485,6.92 sg13_lv_pmos
M$20 \$41 \$14 \$47 \$48 sg13_lv_pmos W=1.4999999999999998 L=0.12999999999999995
* device instance $21 r0 *1 -9.756,4.267 cap_cmim
C$21 \$17 \$41 cap_cmim w=5.77 l=5.77 m=1
* device instance $22 r0 *1 -10.985,12.009 cap_cmim
C$22 \$10 \$17 cap_cmim w=8.16 l=8.16 m=1
* device instance $23 r0 *1 5.365,13.251 cap_cmim
C$23 \$59 \$11 cap_cmim w=8.16 l=8.16 m=1
.ENDS stage_t1
