** sch_path: /foss/designs/week12/IDSM2_t1.sch

.subckt IDSM2_t1 vhi vlo vdda vin dout res clkin
x1 vhi vlo vdda vss vin dout res clkin IDSM2_t1_inner
.ends


.subckt IDSM2_t1_inner vhi vlo vdda vssa vin dout res clkin
*.PININFO clkin:I res:I vin:I vssa:I vdda:I vlo:I vhi:I dd:O
x1 vdda p2 net1 net2 vmid2 dout vssa p1 res vout2 comp_t1
x2 p1e clkin p1 p2 p2e clk_generator_t1
x3 res p1e p1 p2 vhi vdda vin vout1 vssa net2 net3 vlo stage_t1
x4 res p2e p2 p1 vhi vdda vout1 vout2 vssa net1 vmid2 vlo stage_t1
.ends

* expanding   symbol:  /foss/designs/week12/comp_t1.sym # of pins=9
** sym_path: /foss/designs/week12/comp_t1.sym
** sch_path: /foss/designs/week12/comp_t1.sch
.subckt comp_t1 vdda pc d dd vinp dout vssa ps res vinm
*.PININFO pc:I vinp:I ps:I vinm:I vdda:B vssa:B d:O dd:O res:I
M4 vinm_samp ps vinm vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M5 vinm_samp psb vinm vdda sg13_lv_pmos L=0.13u W=6u ng=3 m=1
x3 ps VDD VSS psb sg13g2_inv_1
C1 vinm_samp vssa cap_cmim W=5.77e-6 L=5.77e-6 MF=1
M1 out1m pc vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M2 out1m out1p vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M3 out1p out1m vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M6 out1p pc vdda vdda sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M7 out1m out1p d2p vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M8 d2p pc d1p vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M9 d1p vinp vssa vssa sg13_lv_nmos L=1u W=2u ng=1 m=1
M10 out1p out1m d2m vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M11 d2m pc d1m vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M12 d1m vinm_samp vssa vssa sg13_lv_nmos L=1u W=2u ng=1 m=1
M13 net1 out1p VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M14 net1 net2 VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M15 net2 net1 VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M16 net2 out1m VDD VDD sg13_lv_pmos L=0.13u W=4u ng=1 m=1
M17 net1 net2 net3 VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M18 net2 net1 net4 VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M19 net3 out1p VSS net5 sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M20 net4 out1m VSS VSS sg13_lv_nmos L=0.13u W=2u ng=1 m=1
x1 net2 VDD VSS d sg13g2_buf_2
x2 ps net2 dd net7 net6 VDD VSS sg13g2_dfrbp_2
x4 res VDD VSS net6 sg13g2_inv_1
x5 dd VDD VSS dout sg13g2_inv_2
.ends


* expanding   symbol:  /foss/designs/week12/clk_generator_t1.sym # of pins=5
** sym_path: /foss/designs/week12/clk_generator_t1.sym
** sch_path: /foss/designs/week12/clk_generator_t1.sch
.subckt clk_generator_t1 p1e clkin p1 p2 p2e
*.PININFO clkin:I p2e:O p2:O p1:O p1e:O
x1 clkin VDD VSS clkinb sg13g2_inv_2
x2 clkinbb b2 VDD VSS net11 sg13g2_nand2_2
x3 clkinb VDD VSS clkinbb sg13g2_inv_2
x4 net11 VDD VSS net2 sg13g2_inv_4
x8 b1 clkinb VDD VSS net12 sg13g2_nand2_2
x9 net12 VDD VSS net1 sg13g2_inv_4
x15 net2 VDD VSS net4 sg13g2_inv_4
x16 net1 VDD VSS net3 sg13g2_inv_4
x17 net4 VDD VSS net6 sg13g2_inv_4
x18 net3 VDD VSS net5 sg13g2_inv_4
x19 net6 VDD VSS a1 sg13g2_inv_4
x20 net5 VDD VSS a2 sg13g2_inv_4
x21 a1 VDD VSS p1e sg13g2_inv_4
x22 a2 VDD VSS p2e sg13g2_inv_4
x23 p1e VDD VSS b1 sg13g2_inv_4
x24 p2e VDD VSS b2 sg13g2_inv_4
x25 a1 b1 VDD VSS net7 sg13g2_nand2_2
x26 a2 b2 VDD VSS net8 sg13g2_nand2_2
x5 net7 VDD VSS net9 sg13g2_inv_4
x6 net8 VDD VSS net10 sg13g2_inv_4
x7 net9 VDD VSS p1 sg13g2_inv_8
x10 net10 VDD VSS p2 sg13g2_inv_8
.ends


* expanding   symbol:  /foss/designs/week12/stage_t1.sym # of pins=12
** sym_path: /foss/designs/week12/stage_t1.sym
** sch_path: /foss/designs/week12/stage_t1.sch
.subckt stage_t1 res pse ps pr vhi vdda vin vout vssa d vmid vlo
*.PININFO res:I pse:I ps:I pr:I vhi:B vin:I d:I vlo:B vdda:B vssa:B vout:O vmid:O
x1 ps VDD VSS psb sg13g2_inv_1
x2 d pr VDD VSS gp sg13g2_nand2b_1
M2 vout res vx4 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M3 vx1 gp vhi vdda sg13_lv_pmos L=0.13u W=1.5u ng=1 m=1
M4 vx1 ps vin vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M5 vx1 psb vin vdda sg13_lv_pmos L=0.13u W=6u ng=3 m=1
C2 vx2 vx1 cap_cmim W=5.77e-6 L=5.77e-6 MF=1
x4 pr d VDD VSS gn sg13g2_and2_1
M6 vx1 gn vlo vssa sg13_lv_nmos L=0.13u W=0.5u ng=1 m=1
C3 vx3 vx2 cap_cmim W=8.16e-6 L=8.16e-6 MF=1
M7 vx4 pr vx2 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M8 vx4 ps vx3 vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
C4 vx4 vout cap_cmim W=8.16e-6 L=8.16e-6 MF=1
M9 vx2 pse vmid vssa sg13_lv_nmos L=0.13u W=2u ng=1 m=1
M10 vout vx3 vdda vdda sg13_lv_pmos L=1.5u W=10u ng=4 m=1
M11 vout vx3 vssa vssa sg13_lv_nmos L=1.5u W=2.5u ng=1 m=1
M12 vmid vmid vdda vdda sg13_lv_pmos L=1.5u W=10u ng=4 m=1
M13 vmid vmid vssa vssa sg13_lv_nmos L=1.5u W=2.5u ng=1 m=1
.ends

************************************************************************
*
* Copyright 2023 IHP PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*    https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
************************************************************************

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a21o_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a21o_1 A1 A2 B1 VDD VSS X
*.PININFO A1:I A2:I B1:I X:O VDD:B VSS:B
MN0 net1 A1 net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN1 net2 A2 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN2 net1 B1 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN3 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MP0 net1 B1 net3 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net3 A1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP2 net3 A2 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP3 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a21o_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a21o_2 A1 A2 B1 VDD VSS X
*.PININFO A1:I A2:I B1:I X:O VDD:B VSS:B
MN0 net1 A1 net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN1 net2 A2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 net1 B1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN3 X net1 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MP0 net1 B1 net3 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net3 A1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP2 net3 A2 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP3 X net1 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a21oi_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a21oi_1 A1 A2 B1 VDD VSS Y
*.PININFO A1:I A2:I B1:I Y:O VDD:B VSS:B
MMNB0 Y B1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNA1 sndA1 A2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNA0 Y A1 sndA1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMPB0 Y B1 pndA VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPA1 pndA A2 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPA0 pndA A1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a21oi_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a21oi_2 A1 A2 B1 VDD VSS Y
*.PININFO A1:I A2:I B1:I Y:O VDD:B VSS:B
MMNB0 Y B1 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MMNA1 sndA1 A2 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MMNA0 Y A1 sndA1 VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MMPB0 Y B1 pndA VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MMPA1 pndA A2 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MMPA0 pndA A1 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a221oi_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a221oi_1 A1 A2 B1 B2 C1 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C1:I Y:O VDD:B VSS:B
MMPC0 Y C1 pndB VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPB1 pndB B2 pndA VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPB0 pndB B1 pndA VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPA1 pndA A2 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPA0 pndA A1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMNC0 Y C1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNB1 sndB1 B2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNB0 Y B1 sndB1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNA1 sndA1 A2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNA0 Y A1 sndA1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and2_1 A B VDD VSS X
*.PININFO A:I B:I X:O VDD:B VSS:B
MX0 net4 A net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 X net4 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 net2 B VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 net4 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 VDD net4 X VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 net4 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and2_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and2_2 A B VDD VSS X
*.PININFO A:I B:I X:O VDD:B VSS:B
MX0 net4 A net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 X net4 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX3 net2 B VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 net4 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 VDD net4 X VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX5 net4 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and3_1 A B C VDD VSS X
*.PININFO A:I B:I C:I X:O VDD:B VSS:B
MX0 net3 C VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 X net2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 net2 A net1 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX6 net1 B net3 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX3 X net2 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 net2 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 net2 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 net2 C VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and3_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and3_2 A B C VDD VSS X
*.PININFO A:I B:I C:I X:O VDD:B VSS:B
MX0 net3 C VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX2 X net2 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX5 net2 A net1 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX6 net1 B net3 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX3 X net2 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX1 net2 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 net2 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 net2 C VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and4_1 A B C D VDD VSS X
*.PININFO A:I B:I C:I D:I X:O VDD:B VSS:B
MN4 net17 D VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN3 net16 C net17 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN2 net15 B net16 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN1 net1 A net15 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP4 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP3 net1 D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 net1 C VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP1 net1 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_and4_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_and4_2 A B C D VDD VSS X
*.PININFO A:I B:I C:I D:I X:O VDD:B VSS:B
MN4 net17 D VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN3 net16 C net17 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN2 net15 B net16 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN1 net1 A net15 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP4 X net1 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP3 net1 D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 net1 C VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP1 net1 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_antennanp
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_antennanp A VDD VSS
*.PININFO A:I VDD:B VSS:B
Ddn_1 VSS A dantenna m=1 w=780n l=780n a=608.4f p=3.12u
DD0 A VDD dpantenna m=1 w=1.05u l=1.34u a=1.407p p=4.78u
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_1 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_16
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_16 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=4.44u l=130.00n ng=6
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=11.84u l=130.00n ng=16
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=17.92u l=130.00n ng=16
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=6.72u l=130.00n ng=6
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_2 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=1.48u l=130.00n ng=2
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=2.24u l=130.00n ng=2
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_4 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=2.96u l=130.00n ng=4
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=4.48u l=130.00n ng=4
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=1.68u l=130.00n ng=2
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_buf_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_buf_8 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MN1 net1 A VSS VSS sg13_lv_nmos m=1 w=2.22u l=130.00n ng=3
MN0 X net1 VSS VSS sg13_lv_nmos m=1 w=5.92u l=130.00n ng=8
MP1 X net1 VDD VDD sg13_lv_pmos m=1 w=8.96u l=130.00n ng=8
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=3.36u l=130.00n ng=3
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_decap_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_decap_4 VDD VSS
*.PININFO VDD:B VSS:B
MX1 VSS VDD VSS VSS sg13_lv_nmos m=1 w=420.00n l=1.000u ng=1
MX0 VDD VSS VDD VDD sg13_lv_pmos m=1 w=1.000u l=1.000u ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_decap_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_decap_8 VDD VSS
*.PININFO VDD:B VSS:B
MX1 VSS VDD VSS VSS sg13_lv_nmos m=2 w=420.00n l=1.000u ng=1
MX0 VDD VSS VDD VDD sg13_lv_pmos m=2 w=1.000u l=1.000u ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dfrbp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dfrbp_1 CLK D Q Q_N RESET_B VDD VSS
*.PININFO CLK:I D:I RESET_B:I Q:O Q_N:O VDD:B VSS:B
MN13 net12 net2 VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN14 net5 clkneg net12 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN15 net2 net5 net11 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN16 net11 RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN6 Q_N net5 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 Db D net10 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN1 net10 RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN7 Db clkneg net6 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN8 net6 clkpos net9 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN9 net9 net4 net8 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN10 net8 RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN11 net4 net6 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN2 clkneg CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN12 net4 clkpos net5 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN3 clkpos clkneg VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN4 Q net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN5 net1 net5 VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MP14 net5 clkpos net3 VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP15 net2 net5 VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP16 net2 RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP6 Q_N net5 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP7 Db clkpos net6 VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP0 Db RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP1 Db D VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP8 net7 net4 VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP9 net6 clkneg net7 VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP10 net6 RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP2 clkneg CLK VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP3 clkpos clkneg VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP11 net4 net6 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP12 net4 clkneg net5 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP4 Q net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP13 net3 net2 VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP5 net1 net5 VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dfrbp_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dfrbp_2 CLK D Q Q_N RESET_B VDD VSS
*.PININFO CLK:I D:I RESET_B:I Q:O Q_N:O VDD:B VSS:B
MN13 net12 net2 VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN14 net5 clkneg net12 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN15 net2 net5 net11 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN16 net11 RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN6 Q_N net5 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN0 Db D net10 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN1 net10 RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN7 Db clkneg net6 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN8 net6 clkpos net9 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN9 net9 net4 net8 VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN10 net8 RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN11 net4 net6 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 clkneg CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN12 net4 clkpos net5 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN3 clkpos clkneg VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN4 Q net1 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN5 net1 net5 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MP14 net5 clkpos net3 VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP15 net2 net5 VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP16 net2 RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP6 Q_N net5 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP7 Db clkpos net6 VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP0 Db RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP1 Db D VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP8 net7 net4 VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP9 net6 clkneg net7 VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP10 net6 RESET_B VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP2 clkneg CLK VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP3 clkpos clkneg VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP11 net4 net6 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP12 net4 clkneg net5 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP4 Q net1 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP13 net3 net2 VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MP5 net1 net5 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlhq_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlhq_1 D GATE Q VDD VSS
*.PININFO D:I GATE:I Q:O VDD:B VSS:B
MX17 VDD a_386_326_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX16 a_592_149_ a_685_59_ a_419_392_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX14 a_386_326_ a_592_149_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX12 VDD D a_116_424_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX9 a_562_123_ GATE VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 VDD a_562_123_ a_685_59_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX4 VDD a_386_326_ a_419_392_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX3 a_229_392_ a_562_123_ a_592_149_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n
+ ng=1
MX1 a_229_392_ a_116_424_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX15 a_562_123_ GATE VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX13 VSS a_562_123_ a_685_59_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 a_514_149_ a_562_123_ a_592_149_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX10 VSS a_386_326_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 a_239_85_ a_116_424_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 VSS a_386_326_ a_514_149_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX5 a_386_326_ a_592_149_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 a_592_149_ a_685_59_ a_239_85_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n
+ ng=1
MX0 VSS D a_116_424_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlhr_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlhr_1 D GATE Q Q_N RESET_B VDD VSS
*.PININFO D:I GATE:I RESET_B:I Q:O Q_N:O VDD:B VSS:B
MX0 a_823_98_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 VDD a_823_98_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX15 a_642_392_ a_353_98_ a_753_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX6 a_753_508_ a_823_98_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX10 a_564_392_ a_226_104_ a_642_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n
+ ng=1
MX18 VDD a_27_142_ a_564_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX13 a_27_142_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 VDD GATE a_226_104_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 VDD a_1342_74_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 VDD a_642_392_ a_823_98_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX20 a_353_98_ a_226_104_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX2 a_1342_74_ a_823_98_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX12 a_823_98_ a_642_392_ a_1051_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n
+ ng=1
MX21 a_1051_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX11 a_642_392_ a_226_104_ a_775_124_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX14 a_775_124_ a_823_98_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX7 VSS a_823_98_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 a_571_80_ a_353_98_ a_642_392_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n
+ ng=1
MX23 VSS a_27_142_ a_571_80_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX4 a_27_142_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX19 VSS GATE a_226_104_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 VSS a_1342_74_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 a_353_98_ a_226_104_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 a_1342_74_ a_823_98_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlhrq_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlhrq_1 D GATE Q RESET_B VDD VSS
*.PININFO D:I GATE:I RESET_B:I Q:O VDD:B VSS:B
MX19 a_769_74_ a_817_48_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX14 a_565_74_ a_363_74_ a_643_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n
+ ng=1
MX11 VSS a_817_48_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX10 a_27_424_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX8 a_1045_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 a_817_48_ a_643_74_ a_1045_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n
+ ng=1
MX6 a_643_74_ a_216_424_ a_769_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX4 VSS GATE a_216_424_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 VSS a_27_424_ a_565_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX1 a_363_74_ a_216_424_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 VDD a_643_74_ a_817_48_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX17 VDD a_27_424_ a_568_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX16 a_643_74_ a_363_74_ a_759_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX15 VDD GATE a_216_424_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX13 a_27_424_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX12 a_759_508_ a_817_48_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX9 a_363_74_ a_216_424_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 VDD a_817_48_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_817_48_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX0 a_568_392_ a_216_424_ a_643_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n
+ ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dllr_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dllr_1 D GATE_N Q Q_N RESET_B VDD VSS
*.PININFO D:I GATE_N:I Q:I RESET_B:I Q_N:O VDD:B VSS:B
MX19 VDD a_686_74_ a_889_92_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX17 a_802_508_ a_889_92_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX16 a_27_424_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX11 VDD a_27_424_ a_611_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX10 a_889_92_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX9 a_686_74_ a_231_74_ a_802_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX7 VDD GATE_N a_231_74_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX6 a_1437_112_ a_889_92_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 a_611_392_ a_373_74_ a_686_74_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX3 VDD a_889_92_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 a_373_74_ a_231_74_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 VDD a_1437_112_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX23 VSS a_1437_112_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX22 a_373_74_ a_231_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX21 a_889_92_ a_686_74_ a_1133_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n
+ ng=1
MX20 VSS GATE_N a_231_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 a_1437_112_ a_889_92_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX15 a_27_424_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX14 a_841_118_ a_889_92_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX13 VSS a_27_424_ a_608_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX12 a_686_74_ a_373_74_ a_841_118_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX8 VSS a_889_92_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_608_74_ a_231_74_ a_686_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX0 a_1133_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dllrq_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dllrq_1 D GATE_N Q RESET_B VDD VSS
*.PININFO D:I GATE_N:I RESET_B:I Q:O VDD:B VSS:B
MX18 a_357_392_ a_232_98_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX17 VSS a_897_406_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 a_654_392_ a_357_392_ a_854_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX14 VSS a_27_136_ a_681_74_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX12 a_681_74_ a_232_98_ a_654_392_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n
+ ng=1
MX9 a_27_136_ D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX6 a_1139_74_ RESET_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 a_854_74_ a_897_406_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX3 a_897_406_ a_654_392_ a_1139_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n
+ ng=1
MX1 VSS GATE_N a_232_98_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX19 VDD GATE_N a_232_98_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX15 a_897_406_ RESET_B VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX13 a_654_392_ a_232_98_ a_793_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX11 a_793_508_ a_897_406_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX10 VDD a_897_406_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX8 a_27_136_ D VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 VDD a_27_136_ a_570_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 VDD a_654_392_ a_897_406_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX2 a_570_392_ a_357_392_ a_654_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n
+ ng=1
MX0 a_357_392_ a_232_98_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlygate4sd1_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlygate4sd1_1 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MP3 X net3 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP2 net3 net2 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net2 net1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MN3 X net3 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 net3 net2 VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN1 net2 net1 VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN0 net1 A VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlygate4sd2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlygate4sd2_1 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MP3 X net3 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP2 net3 net2 VDD VDD sg13_lv_pmos m=1 w=1.000u l=250.00n ng=1
MP1 net2 net1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=250.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MN3 X net3 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 net3 net2 VSS VSS sg13_lv_nmos m=1 w=420.00n l=180.00n ng=1
MN1 net2 net1 VSS VSS sg13_lv_nmos m=1 w=420.00n l=180.00n ng=1
MN0 net1 A VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_dlygate4sd3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_dlygate4sd3_1 A VDD VSS X
*.PININFO A:I X:O VDD:B VSS:B
MP3 X net3 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP2 net3 net2 VDD VDD sg13_lv_pmos m=1 w=1.000u l=500.0n ng=1
MP1 net2 net1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=500.0n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MN3 X net3 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 net3 net2 VSS VSS sg13_lv_nmos m=1 w=420.00n l=500.0n ng=1
MN1 net2 net1 VSS VSS sg13_lv_nmos m=1 w=420.00n l=500.0n ng=1
MN0 net1 A VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_ebufn_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_ebufn_2 A TE_B VDD VSS Z
*.PININFO A:I TE_B:I Z:O VDD:B VSS:B
MN3 net4 net3 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN2 Z net1 net4 VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN1 net3 TE_B VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN0 net1 A VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MP3 net2 TE_B VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP2 Z net1 net2 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP1 net3 TE_B VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_ebufn_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_ebufn_4 A TE_B VDD VSS Z
*.PININFO A:I TE_B:I Z:O VDD:B VSS:B
MN0 net23 A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN1 net21 TE_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 Z net23 net22 VSS sg13_lv_nmos m=4 w=740.00n l=130.00n ng=1
MN3 net22 net21 VSS VSS sg13_lv_nmos m=4 w=740.00n l=130.00n ng=1
MP0 net23 A VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP1 net21 TE_B VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP2 Z net23 net24 VDD sg13_lv_pmos m=4 w=1.12u l=130.00n ng=1
MP3 net24 TE_B VDD VDD sg13_lv_pmos m=4 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_ebufn_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_ebufn_8 A TE_B VDD VSS Z
*.PININFO A:I TE_B:I Z:O VDD:B VSS:B
MN3 net23 net22 VSS VSS sg13_lv_nmos m=8 w=740.00n l=130.00n ng=1
MN2 Z net21 net23 VSS sg13_lv_nmos m=8 w=740.00n l=130.00n ng=1
MN1 net22 TE_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 net21 A VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MP3 net24 TE_B VDD VDD sg13_lv_pmos m=8 w=1.12u l=130.00n ng=1
MP2 Z net21 net24 VDD sg13_lv_pmos m=8 w=1.12u l=130.00n ng=1
MP1 net22 TE_B VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP0 net21 A VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_einvn_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_einvn_2 A TE_B VDD VSS Z
*.PININFO A:I TE_B:I Z:O VDD:B VSS:B
MN2 TE TE_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MN1 net1 TE VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN0 Z A net1 VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MP2 TE TE_B VDD VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MP1 net2 TE_B VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP0 Z A net2 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_einvn_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_einvn_4 A TE_B VDD VSS Z
*.PININFO A:I TE_B:I Z:O VDD:B VSS:B
MN1 net16 TE VSS VSS sg13_lv_nmos m=4 w=740.00n l=130.00n ng=1
MN2 TE TE_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 Z A net16 VSS sg13_lv_nmos m=4 w=740.00n l=130.00n ng=1
MP2 TE TE_B VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP1 net17 TE_B VDD VDD sg13_lv_pmos m=4 w=1.12u l=130.00n ng=1
MP0 Z A net17 VDD sg13_lv_pmos m=4 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_einvn_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_einvn_8 A TE_B VDD VSS Z
*.PININFO A:I TE_B:I Z:O VDD:B VSS:B
MN0 Z A net29 VSS sg13_lv_nmos m=8 w=740.00n l=130.00n ng=1
MN2 TE TE_B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN1 net29 TE VSS VSS sg13_lv_nmos m=8 w=740.00n l=130.00n ng=1
MP1 net28 TE_B VDD VDD sg13_lv_pmos m=8 w=1.12u l=130.00n ng=1
MP0 Z A net28 VDD sg13_lv_pmos m=8 w=1.12u l=130.00n ng=1
MP2 TE TE_B VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_1 A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MX1 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX0 Y A VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_16
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_16 A VSS VDD Y
*.PININFO A:I Y:O VDD:B VSS:B
MX1 Y A VSS VSS sg13_lv_nmos m=16 w=740.00n l=130.00n ng=1
MX0 Y A VDD VDD sg13_lv_pmos m=16 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_2 A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MX1 Y A VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX0 Y A VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_4
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_4 A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MP0 Y A VDD VDD sg13_lv_pmos m=4 w=1.12u l=130.00n ng=1
MN0 Y A VSS VSS sg13_lv_nmos m=4 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_inv_8
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_inv_8 A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MX1 Y A VSS VSS sg13_lv_nmos m=8 w=740.00n l=130.00n ng=1
MX0 Y A VDD VDD sg13_lv_pmos m=8 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_lgcp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_lgcp_1 CLK GATE GCLK VDD VSS
*.PININFO CLK:I GATE:I GCLK:O VDD:B VSS:B
MX15 CLKBB CLKB VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX14 a_83_260_ CLKBB a_258_392_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX12 int_GATE a_83_260_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX11 a_258_392_ GATE VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX9 a_987_393_ int_GATE VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 GCLK a_987_393_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 a_83_260_ CLKB a_484_508_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX4 CLKB CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 a_987_393_ CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX2 a_484_508_ int_GATE VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX19 GCLK a_987_393_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 a_987_393_ int_GATE a_984_125_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n
+ ng=1
MX17 int_GATE a_83_260_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX16 CLKBB CLKB VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX13 a_477_124_ int_GATE VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 a_267_80_ GATE VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 a_83_260_ CLKBB a_477_124_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX6 CLKB CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 a_984_125_ CLK VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX0 a_83_260_ CLKB a_267_80_ VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_mux2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_mux2_1 A0 A1 S VDD VSS X
*.PININFO A0:I A1:I S:I X:O VDD:B VSS:B
MP0 net4 S VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP4 X net6 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP3 net6 A1 net5 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP5 Sb S VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 net5 Sb VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net6 A0 net4 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MN4 net3 S VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN1 net1 Sb VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN6 X net6 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN5 Sb S VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 net6 A1 net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 net6 A0 net1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_mux2_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_mux2_2 A0 A1 S VDD VSS X
*.PININFO A0:I A1:I S:I X:O VDD:B VSS:B
MP0 net4 S VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP4 X net6 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP3 net6 A1 net5 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP5 Sb S VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 net5 Sb VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net6 A0 net4 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MN4 net3 S VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN1 net1 Sb VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN6 X net6 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN5 Sb S VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 net6 A1 net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 net6 A0 net1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_mux4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_mux4_1 A0 A1 A2 A3 S0 S1 VDD VSS X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I X:O VDD:B VSS:B
MN12 X Xb VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN18 low S0b net7 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN17 net7 A0 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN19 low S1b Xb VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN10 high S1 Xb VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN9 net4 A3 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN8 high S0 net4 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN14 net6 A2 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN13 high S0b net6 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN16 net2 A1 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN15 low S0 net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN1 S1b S1 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN0 S0b S0 VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MP19 low S1 Xb VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP11 high S1b Xb VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP10 X Xb VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP9 high S0b net3 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP8 net3 A3 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP14 high S0 net5 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP13 net5 A2 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP18 net8 A0 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP17 low S0 net8 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 S1b S1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP0 S0b S0 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP16 low S0b net1 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP15 net1 A1 VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand2_1 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MP1 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MP0 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MN1 net1 B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 Y A net1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand2_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand2_2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MP1 Y B VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MP0 Y A VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MN1 net1 B VSS VSS sg13_lv_nmos m=2 w=720.00n l=130.00n ng=1
MN0 Y A net1 VSS sg13_lv_nmos m=2 w=720.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand2b_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand2b_1 A_N B VDD VSS Y
*.PININFO A_N:I B:I Y:O VDD:B VSS:B
MX0 Y a_27_112_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 a_27_112_ A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y a_27_112_ net1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_27_112_ A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX5 net1 B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand2b_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand2b_2 A_N B VDD VSS Y
*.PININFO A_N:I B:I Y:O VDD:B VSS:B
MX0 Y A VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX1 A A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 Y B VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX2 Y A net1 VSS sg13_lv_nmos m=2 w=720.00n l=130.00n ng=1
MX4 A A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX5 net1 B VSS VSS sg13_lv_nmos m=2 w=720.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand3_1 A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MX1 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 Y C VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net2 B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 net3 C VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 Y A net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand3b_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand3b_1 A_N B C VDD VSS Y
*.PININFO A_N:I B:I C:I Y:O VDD:B VSS:B
MX0 net1 A_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 Y net1 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 Y C VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net2 B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 net3 C VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX5 net1 A_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 Y net1 net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nand4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nand4_1 A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MP0 Y D VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 Y C VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net2 B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 net3 C net5 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX7 Y A net2 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN0 net5 D VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor2_1 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MX0 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 Y B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX1 net1 A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B net1 VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor2_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor2_2 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MX0 Y A VSS VSS sg13_lv_nmos m=1 w=1.48u l=130.00n ng=2
MX3 Y B VSS VSS sg13_lv_nmos m=1 w=1.48u l=130.00n ng=2
MX1 net1 A VDD VDD sg13_lv_pmos m=1 w=2.24u l=130.00n ng=2
MX2 Y B net1 VDD sg13_lv_pmos m=1 w=2.24u l=130.00n ng=2
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor2b_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor2b_1 A B_N VDD VSS Y
*.PININFO A:I B_N:I Y:O VDD:B VSS:B
MN0 B B_N VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX0 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 Y B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MP0 B B_N VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX1 net1 A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX2 Y B net1 VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor2b_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor2b_2 A B_N VDD VSS Y
*.PININFO A:I B_N:I Y:O VDD:B VSS:B
MN0 B B_N VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX0 Y A VSS VSS sg13_lv_nmos m=2 w=720.00n l=130.00n ng=1
MX3 Y B VSS VSS sg13_lv_nmos m=2 w=720.00n l=130.00n ng=1
MP0 B B_N VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX1 net1 A VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX2 Y B net1 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor3_1 A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MX3 net1 C Y VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MX0 net2 B net1 VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MX2 VDD A net2 VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MX4 Y A VSS VSS sg13_lv_nmos m=1 w=770.00n l=130.00n ng=1
MX1 Y B VSS VSS sg13_lv_nmos m=1 w=770.00n l=130.00n ng=1
MX5 Y C VSS VSS sg13_lv_nmos m=1 w=770.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor3_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor3_2 A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MX3 net1 C Y VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX0 net2 B net1 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX2 VDD A net2 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX4 Y A VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX1 Y B VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX5 Y C VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor4_1 A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MX0 net3 A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 net2 B net3 VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX6 net1 C net2 VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 Y D net1 VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX1 Y A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX2 Y D VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX3 Y B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 Y C VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_nor4_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_nor4_2 A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MX0 net3 A VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX5 net2 B net3 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX6 net1 C net2 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX7 Y D net1 VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX1 Y A VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX2 Y D VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX3 Y B VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX4 Y C VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_o21ai_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_o21ai_1 A1 A2 B1 VDD VSS Y
*.PININFO A1:I A2:I B1:I Y:O VDD:B VSS:B
MP2 net14 A1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=150.00n ng=1
MP1 Y A2 net14 VDD sg13_lv_pmos m=1 w=1.12u l=150.00n ng=1
MP0 Y B1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=150.00n ng=1
MN2 net1 A2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=150.00n ng=1
MN3 net1 A1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=150.00n ng=1
MN0 Y B1 net1 VSS sg13_lv_nmos m=1 w=740.00n l=150.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or2_1 A B VDD VSS X
*.PININFO A:I B:I X:O VDD:B VSS:B
MP0 net2 B net3 VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP1 net3 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 X net2 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MN0 net2 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN1 net2 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 X net2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or2_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or2_2 A B VDD VSS X
*.PININFO A:I B:I X:O VDD:B VSS:B
MP0 net2 B net3 VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP1 net3 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP2 X net2 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MN0 net2 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN1 net2 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 X net2 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or3_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or3_1 A B C VDD VSS X
*.PININFO A:I B:I C:I X:O VDD:B VSS:B
MX0 net1 C VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 net1 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX2 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX3 net9 B net12 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 net12 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX5 net1 C net9 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or3_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or3_2 A B C VDD VSS X
*.PININFO A:I B:I C:I X:O VDD:B VSS:B
MX0 net1 C VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 X net1 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MX6 net1 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX7 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX2 X net1 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
MX3 net9 B net12 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX4 net12 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX5 net1 C net9 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or4_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or4_1 A B C D VDD VSS X
*.PININFO A:I B:I C:I D:I X:O VDD:B VSS:B
MN4 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN3 net1 D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 net1 C VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN1 net1 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN0 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MP4 net4 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP3 net3 B net4 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP2 net2 C net3 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net1 D net2 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP0 X net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_or4_2
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_or4_2 A B C D VDD VSS X
*.PININFO A:I B:I C:I D:I X:O VDD:B VSS:B
MN4 X net1 VSS VSS sg13_lv_nmos m=2 w=740.00n l=130.00n ng=1
MN3 net1 D VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN2 net1 C VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN1 net1 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MN0 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MP4 net4 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP3 net3 B net4 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP2 net2 C net3 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP1 net1 D net2 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MP0 X net1 VDD VDD sg13_lv_pmos m=2 w=1.12u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_sdfbbp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_sdfbbp_1 CLK D Q Q_N RESET_B SCD SCE SET_B VDD VSS
*.PININFO CLK:I D:I RESET_B:I SCD:I SCE:I SET_B:I Q:O Q_N:O VDD:B VSS:B
MX46 a_1625_93_ RESET_B VDD VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX45 a_2037_442_ a_1878_420_ a_2384_392_ VDD sg13_lv_pmos m=1 w=1.000u
+ l=130.00n ng=1
MX44 VDD SET_B a_2037_442_ VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX41 VDD a_622_98_ a_877_98_ VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX39 VDD SCE a_341_93_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX38 a_218_464_ D a_197_119_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX33 a_1092_96_ a_622_98_ a_1221_419_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX28 a_1221_419_ a_1250_231_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX27 VDD SCE a_218_464_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX26 VDD a_2037_442_ Q_N VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX24 VDD a_1250_231_ a_1766_379_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX19 a_2384_392_ a_1625_93_ VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX17 VDD SET_B a_1250_231_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX16 a_27_464_ SCD VDD VDD sg13_lv_pmos m=1 w=640.00n l=130.00n ng=1
MX15 a_622_98_ CLK VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX14 a_1250_231_ a_1092_96_ a_1580_379_ VDD sg13_lv_pmos m=1 w=840.00n
+ l=130.00n ng=1
MX11 a_197_119_ a_877_98_ a_1092_96_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n
+ ng=1
MX9 a_197_119_ a_341_93_ a_27_464_ VDD sg13_lv_pmos m=1 w=640.00n l=130.00n
+ ng=1
MX8 a_2881_74_ a_2037_442_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX7 a_1580_379_ a_1625_93_ VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX6 a_1986_504_ a_2037_442_ VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX5 a_1878_420_ a_877_98_ a_1986_504_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n
+ ng=1
MX4 a_1766_379_ a_622_98_ a_1878_420_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n
+ ng=1
MX3 VDD a_2881_74_ Q VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX47 a_2271_74_ a_1878_420_ a_2037_442_ VSS sg13_lv_nmos m=1 w=740.00n
+ l=130.00n ng=1
MX43 a_197_119_ a_622_98_ a_1092_96_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX42 a_299_119_ a_341_93_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX40 VSS a_622_98_ a_877_98_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX37 a_1625_93_ RESET_B VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX36 a_2061_74_ a_2037_442_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX35 a_1418_125_ a_1092_96_ a_1250_231_ VSS sg13_lv_nmos m=1 w=550.00n
+ l=130.00n ng=1
MX34 VSS SCE a_341_93_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX32 VSS SET_B a_1418_125_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX31 a_1192_96_ a_1250_231_ VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX30 a_119_119_ SCE a_197_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX29 VSS SET_B a_2271_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX25 a_1092_96_ a_877_98_ a_1192_96_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX23 a_197_119_ D a_299_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX22 a_2881_74_ a_2037_442_ VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX21 a_1878_420_ a_622_98_ a_2061_74_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n
+ ng=1
MX20 VSS a_2881_74_ Q VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX18 VSS a_1250_231_ a_1880_119_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX13 a_622_98_ CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX12 VSS SCD a_119_119_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 a_1880_119_ a_877_98_ a_1878_420_ VSS sg13_lv_nmos m=1 w=550.00n
+ l=130.00n ng=1
MX2 a_1250_231_ a_1625_93_ a_1418_125_ VSS sg13_lv_nmos m=1 w=550.00n
+ l=130.00n ng=1
MX1 VSS a_2037_442_ Q_N VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX0 a_2037_442_ a_1625_93_ a_2271_74_ VSS sg13_lv_nmos m=1 w=740.00n l=130.00n
+ ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_sighold
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_sighold SH VDD VSS
*.PININFO SH:B VDD:B VSS:B
MN0 net1 SH VSS VSS sg13_lv_nmos m=1 w=300.0n l=130.00n ng=1
MN1 SH net1 VSS VSS sg13_lv_nmos m=1 w=300.0n l=700.0n ng=1
MP0 net1 SH VDD VDD sg13_lv_pmos m=1 w=450.00n l=130.00n ng=1
MP1 SH net1 VDD VDD sg13_lv_pmos m=1 w=300.0n l=700.0n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_slgcp_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_slgcp_1 CLK GATE GCLK SCE VDD VSS
*.PININFO CLK:I GATE:I SCE:I GCLK:O VDD:B VSS:B
MX19 GCLK a_1238_94_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX18 a_114_112_ CLKbb a_566_74_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX16 CLKbb CLKb VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX14 a_1238_94_ int_GATE VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX13 a_116_424_ SCE VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX11 a_566_74_ CLKb a_722_492_ VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX9 int_GATE a_566_74_ VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 CLKb CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX5 a_1238_94_ CLK VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX3 a_722_492_ int_GATE VDD VDD sg13_lv_pmos m=1 w=420.00n l=130.00n ng=1
MX2 a_114_112_ GATE a_116_424_ VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MX21 int_GATE a_566_74_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX20 net2 CLK VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX17 a_114_112_ SCE VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX15 a_566_74_ CLKb a_114_112_ VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX12 a_667_80_ int_GATE VSS VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
MX10 a_1238_94_ int_GATE net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MX8 GCLK a_1238_94_ VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 CLKbb CLKb VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX4 a_114_112_ GATE VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 CLKb CLK VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX0 a_566_74_ CLKbb a_667_80_ VSS sg13_lv_nmos m=1 w=420.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_tiehi
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_tiehi L_HI VDD VSS
*.PININFO L_HI:O VDD:B VSS:B
MMN2 net3 net2 VSS VSS sg13_lv_nmos m=1 w=795.00n l=130.00n ng=1
MMN1 net1 net1 VSS VSS sg13_lv_nmos m=1 w=300n l=130.00n ng=1
MMP2 L_HI net3 VDD VDD sg13_lv_pmos m=1 w=1.155u l=130.00n ng=1
MMP1 net2 net1 VDD VDD sg13_lv_pmos m=1 w=660.0n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_tielo
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_tielo L_LO VDD VSS
*.PININFO L_LO:O VDD:B VSS:B
MMN1 net3 net2 VSS VSS sg13_lv_nmos m=1 w=385.00n l=130.00n ng=1
MMN2 L_LO net1 VSS VSS sg13_lv_nmos m=1 w=880.0n l=130.00n ng=1
MMP1 net2 net2 VDD VDD sg13_lv_pmos m=1 w=300n l=130.00n ng=1
MMP2 net1 net3 VDD VDD sg13_lv_pmos m=1 w=1.045u l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_xnor2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_xnor2_1 A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MP9 Y net1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP8 Y B net4 VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP7 net4 A VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MP1 net1 B VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MP0 net1 A VDD VDD sg13_lv_pmos m=1 w=840.00n l=130.00n ng=1
MN4 Y net1 net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN6 net2 A VSS VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN5 net1 B net2 VSS sg13_lv_nmos m=1 w=640.00n l=130.00n ng=1
MN3 net3 B VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MN2 net3 A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_xor2_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_xor2_1 A B VDD VSS X
*.PININFO A:I B:I X:O VDD:B VSS:B
MX0 net1 A VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX4 X B net3 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX6 X net1 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX8 net3 A VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MX9 net1 B VSS VSS sg13_lv_nmos m=1 w=550.00n l=130.00n ng=1
MX1 net6 A VDD VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX2 net1 B net6 VDD sg13_lv_pmos m=1 w=1.000u l=130.00n ng=1
MX3 net5 A VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX5 net5 B VDD VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
MX7 X net1 net5 VDD sg13_lv_pmos m=1 w=1.12e-06 l=130.00n ng=1
.ENDS

************************************************************************
* Library Name: sg13g2_stdcell
* Cell Name:    sg13g2_a22oi_1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_a22oi_1 A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MN3 net1 B2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNB0 Y B1 net1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNA1 sndA1 A2 VSS VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MMNA0 Y A1 sndA1 VSS sg13_lv_nmos m=1 w=740.00n l=130.00n ng=1
MP3 Y B1 pndA VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPB0 Y B2 pndA VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPA1 pndA A2 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
MMPA0 pndA A1 VDD VDD sg13_lv_pmos m=1 w=1.12u l=130.00n ng=1
.ENDS

.GLOBAL VDD
.GLOBAL VSS
.end
