* Extracted by KLayout with SG13G2 LVS runset on : 06/05/2024 21:09

* cell stage_t1
* pin d
* pin pr
* pin ps
* pin VMID
* pin Vout
* pin VDD
* pin VLO
* pin Vin
* pin VDDA
* pin VHI
* pin VSS
.SUBCKT stage_t1 d pr ps VMID Vout VDD VLO Vin VDDA VHI VSS
* device instance $1 r0 *1 -8.975,-0.35 sg13_lv_nmos
M$1 VSS ps \$12 VSS sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $2 r0 *1 -7.89,-0.25 sg13_lv_nmos
M$2 VSS d \$13 VSS sg13_lv_nmos W=0.5499999999999999 L=0.12999999999999995
* device instance $3 r0 *1 -7.04,-0.345 sg13_lv_nmos
M$3 VSS pr \$22 VSS sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $4 r0 *1 -6.73,-0.345 sg13_lv_nmos
M$4 \$22 \$13 \$14 VSS sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $5 r0 *1 -5.415,-0.18 sg13_lv_nmos
M$5 \$17 pr \$24 VSS sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $6 r0 *1 -4.905,-0.18 sg13_lv_nmos
M$6 VSS d \$24 VSS sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $7 r0 *1 -4.395,-0.23 sg13_lv_nmos
M$7 VSS \$17 \$15 VSS sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $8 r0 *1 12.911,0.09 sg13_lv_nmos
M$8 \$10 \$27 \$16 VSS sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $9 r0 *1 13.42,0.09 sg13_lv_nmos
M$9 \$16 \$28 Vout VSS sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $10 r0 *1 8.511,0.11 sg13_lv_nmos
M$10 VMID \$19 \$18 VSS sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $11 r0 *1 9.02,0.11 sg13_lv_nmos
M$11 \$18 \$20 \$16 VSS sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $12 r0 *1 13.23,2.985 sg13_lv_nmos
M$12 VSS \$10 Vout VSS sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $13 r0 *1 8.855,3 sg13_lv_nmos
M$13 VSS VMID VMID VSS sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $14 r0 *1 0.414,3.383 sg13_lv_nmos
M$14 VLO \$15 \$38 VSS sg13_lv_nmos W=0.4999999999999999 L=0.12999999999999998
* device instance $15 r0 *1 2.832,3.445 sg13_lv_nmos
M$15 \$38 ps Vin VSS sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $16 r0 *1 -7.89,1.175 sg13_lv_pmos
M$16 \$13 d VDD VDD sg13_lv_pmos W=0.8399999999999999 L=0.12999999999999995
* device instance $17 r0 *1 -7.35,1.315 sg13_lv_pmos
M$17 VDD pr \$14 VDD sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $18 r0 *1 -6.84,1.315 sg13_lv_pmos
M$18 \$14 \$13 VDD VDD sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $19 r0 *1 -5.415,1.46 sg13_lv_pmos
M$19 VDD pr \$17 VDD sg13_lv_pmos W=0.8399999999999999 L=0.12999999999999995
* device instance $20 r0 *1 -4.905,1.46 sg13_lv_pmos
M$20 VDD d \$17 VDD sg13_lv_pmos W=0.8399999999999999 L=0.12999999999999995
* device instance $21 r0 *1 -4.395,1.32 sg13_lv_pmos
M$21 VDD \$17 \$15 VDD sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $22 r0 *1 -8.965,1.325 sg13_lv_pmos
M$22 VDD ps \$12 VDD sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $23 r0 *1 13.236,5.995 sg13_lv_pmos
M$23 \$44 \$10 VDDA VDDA sg13_lv_pmos W=2.4999999999999996 L=1.4999999999999996
* device instance $24 r0 *1 13.236,7.875 sg13_lv_pmos
M$24 VDDA \$10 Vout VDDA sg13_lv_pmos W=7.499999999999998 L=1.4999999999999996
* device instance $27 r0 *1 8.866,6.01 sg13_lv_pmos
M$27 VMID VMID VDDA VDDA sg13_lv_pmos W=9.999999999999998 L=1.4999999999999996
* device instance $31 r0 *1 0.818,6.277 sg13_lv_pmos
M$31 \$38 \$12 Vin VDDA sg13_lv_pmos W=5.999999999999998 L=0.12999999999999998
* device instance $34 r0 *1 3.485,6.92 sg13_lv_pmos
M$34 \$38 \$14 VHI VDDA sg13_lv_pmos W=1.4999999999999998 L=0.12999999999999995
* device instance $35 r0 *1 -9.737,4.316 cap_cmim
C$35 \$18 \$38 cap_cmim w=5.77 l=5.77 m=1
* device instance $36 r0 *1 -10.985,12.009 cap_cmim
C$36 \$10 \$18 cap_cmim w=8.16 l=8.16 m=1
* device instance $37 r0 *1 5.365,13.251 cap_cmim
C$37 \$59 Vout cap_cmim w=8.16 l=8.16 m=1
.ENDS stage_t1
