* Extracted by KLayout with SG13G2 LVS runset on : 06/05/2024 00:44

* cell stage_t1
* pin sub!
.SUBCKT stage_t1 sub!
* device instance $1 r0 *1 -8.975,-0.35 sg13_lv_nmos
M$1 sub! \$5 \$13 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $2 r0 *1 -7.89,-0.25 sg13_lv_nmos
M$2 sub! \$1 \$14 sub! sg13_lv_nmos W=0.5499999999999999 L=0.12999999999999995
* device instance $3 r0 *1 -7.04,-0.345 sg13_lv_nmos
M$3 sub! \$2 \$20 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $4 r0 *1 -6.73,-0.345 sg13_lv_nmos
M$4 \$20 \$14 \$15 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $5 r0 *1 -5.415,-0.18 sg13_lv_nmos
M$5 \$16 \$2 \$22 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $6 r0 *1 -4.905,-0.18 sg13_lv_nmos
M$6 sub! \$1 \$22 sub! sg13_lv_nmos W=0.6399999999999999 L=0.12999999999999995
* device instance $7 r0 *1 -4.395,-0.23 sg13_lv_nmos
M$7 sub! \$16 \$17 sub! sg13_lv_nmos W=0.7399999999999999 L=0.12999999999999995
* device instance $8 r0 *1 12.911,0.09 sg13_lv_nmos
M$8 \$11 \$27 \$10 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $9 r0 *1 13.42,0.09 sg13_lv_nmos
M$9 \$10 \$28 \$12 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $10 r0 *1 8.511,0.11 sg13_lv_nmos
M$10 \$9 \$24 \$18 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $11 r0 *1 9.02,0.11 sg13_lv_nmos
M$11 \$18 \$25 \$10 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $12 r0 *1 13.23,2.985 sg13_lv_nmos
M$12 sub! \$11 \$12 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $13 r0 *1 8.855,3 sg13_lv_nmos
M$13 sub! \$9 \$42 sub! sg13_lv_nmos W=2.4999999999999996 L=1.4999999999999996
* device instance $14 r0 *1 0.414,3.383 sg13_lv_nmos
M$14 \$35 \$17 \$38 sub! sg13_lv_nmos W=0.4999999999999999 L=0.12999999999999998
* device instance $15 r0 *1 2.832,3.445 sg13_lv_nmos
M$15 \$41 \$5 \$39 sub! sg13_lv_nmos W=1.9999999999999996 L=0.12999999999999998
* device instance $16 r0 *1 -7.89,1.175 sg13_lv_pmos
M$16 \$14 \$1 \$26 \$26 sg13_lv_pmos W=0.8399999999999999 L=0.12999999999999995
* device instance $17 r0 *1 -7.35,1.315 sg13_lv_pmos
M$17 \$26 \$2 \$15 \$26 sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $18 r0 *1 -6.84,1.315 sg13_lv_pmos
M$18 \$15 \$14 \$26 \$26 sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $19 r0 *1 -5.415,1.46 sg13_lv_pmos
M$19 \$26 \$2 \$16 \$26 sg13_lv_pmos W=0.8399999999999999 L=0.12999999999999995
* device instance $20 r0 *1 -4.905,1.46 sg13_lv_pmos
M$20 \$26 \$1 \$16 \$26 sg13_lv_pmos W=0.8399999999999999 L=0.12999999999999995
* device instance $21 r0 *1 -4.395,1.32 sg13_lv_pmos
M$21 \$26 \$16 \$17 \$26 sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $22 r0 *1 -8.965,1.325 sg13_lv_pmos
M$22 \$26 \$5 \$13 \$26 sg13_lv_pmos W=1.1199999999999999 L=0.12999999999999995
* device instance $23 r0 *1 13.236,5.995 sg13_lv_pmos
M$23 \$46 \$11 \$47 \$47 sg13_lv_pmos W=2.4999999999999996 L=1.4999999999999996
* device instance $24 r0 *1 13.236,7.875 sg13_lv_pmos
M$24 \$47 \$11 \$12 \$47 sg13_lv_pmos W=7.499999999999998 L=1.4999999999999996
* device instance $27 r0 *1 8.866,6.01 sg13_lv_pmos
M$27 \$42 \$9 \$47 \$47 sg13_lv_pmos W=9.999999999999998 L=1.4999999999999996
* device instance $31 r0 *1 0.818,6.277 sg13_lv_pmos
M$31 \$41 \$13 \$39 \$47 sg13_lv_pmos W=5.999999999999998 L=0.12999999999999998
* device instance $34 r0 *1 3.485,6.92 sg13_lv_pmos
M$34 \$41 \$15 \$49 \$47 sg13_lv_pmos W=1.4999999999999998 L=0.12999999999999995
* device instance $35 r0 *1 5.365,13.251 cap_cmim
C$35 \$59 \$60 cap_cmim w=6.99 l=6.99 m=1
.ENDS stage_t1
